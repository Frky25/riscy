
// Copyright (c) 2017 Massachusetts Institute of Technology

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

`include "ProcConfig.bsv"

import CoreStates::*;

import GetPut::*;

import Abstraction::*;
import RVExec::*;
import RVTypes::*;

import RVAlu::*;
import RVControl::*;
import RVMemory::*;
`ifdef CONFIG_M
import RVMulDiv::*;
`endif

import Btb::*;

interface ExecStage;
endinterface

typedef struct {
    Reg#(Maybe#(FetchState)) fs;
    Reg#(Maybe#(RegFetchState)) rs;
    Reg#(Maybe#(ExecuteState)) es;
    Reg#(Maybe#(WriteBackState)) ws;
    Put#(RVDMemReq) dmemreq;
`ifdef CONFIG_M
    MulDivExec mulDiv;
`endif
    NextAddrPred btb;
} ExecRegs;

module mkExecStage#(ExecRegs er)(ExecStage);

    let dmemreq = er.dmemreq;
`ifdef CONFIG_M
    let mulDiv = er.mulDiv;
`endif
    let btb = er.btb;

    rule doExecute(er.es matches tagged Valid .executeState
                    &&& er.ws == tagged Invalid);
        // get and clear the execute state
        let poisoned = executeState.poisoned;
        let pc = executeState.pc;
        let ppc = executeState.ppc;
        Maybe#(TrapCause) trap = executeState.trap;
        let dInst = executeState.dInst;
        let rVal1 = executeState.rVal1;
        let rVal2 = executeState.rVal2;
        Data data = ?;
        Addr addr = ?;
        er.es <= tagged Invalid;
        
        if (!poisoned) begin
            // execute instruction
            let execResult = basicExec(dInst, rVal1, rVal2, pc);
            data = execResult.data;
            addr = execResult.addr;
            let nextPc = execResult.nextPc;

            //$display("[Exec] pc: 0x%0x, dInst: ", pc, fshow(dInst));
            // check for next address alignment
            if (nextPc[1:0] != 0 && trap == tagged Invalid) begin
                trap = tagged Valid (tagged Exception InstAddrMisaligned);
            end

`ifdef CONFIG_M
            if (dInst.execFunc matches tagged MulDiv .mulDivInst &&& trap == tagged Invalid) begin
                mulDiv.exec(mulDivInst, rVal1, rVal2);
            end
`endif

            if (dInst.execFunc matches tagged Mem .memInst &&& trap == tagged Invalid) begin
                // check allignment
                Bool aligned = (case (memInst.size)
                                    B: True;
                                    H: (execResult.addr[0] == 0);
                                    W: (execResult.addr[1:0] == 0);
                                    D: (execResult.addr[2:0] == 0);
                                endcase);
                if (aligned) begin
                    // send the request to the memory
                    dmemreq.put( RVDMemReq {
                        op: dInst.execFunc.Mem.op,
                        size: dInst.execFunc.Mem.size,
                        isUnsigned: dInst.execFunc.Mem.isUnsigned,
                        addr: zeroExtend(addr),
                        data: data } );
                end else begin
                    // misaligned address exception
                    if ((memInst.op == tagged Mem Ld) || (memInst.op == tagged Mem Lr)) begin
                        trap = tagged Valid (tagged Exception LoadAddrMisaligned);
                    end else begin
                        trap = tagged Valid (tagged Exception StoreAddrMisaligned);
                    end
                end
            end

            // update next pc for fetch stage if no trap and misprediction
            if (trap == tagged Invalid) begin
                if(nextPc != ppc) begin //misprediction
                    //kill invalid instruction in reg fetch
                    if(er.rs matches tagged Valid .validRegFetchState) begin
                        let vrs = validRegFetchState;
                        vrs.poisoned = True;
                        er.rs <= tagged Valid vrs;
                    end
                    //update BTB
                    btb.update(pc, nextPc, pc+4 != nextPc);
                    //correct pc    
                    er.fs <= tagged Valid FetchState{ pc: nextPc };
                end
            end
        end
        
        //always store things for next stage because of bookkeeping
        er.ws <= tagged Valid WriteBackState{
                                            poisoned: poisoned,
                                            pc: pc,
                                            trap: trap,
                                            dInst: dInst,
                                            addr: addr,
                                            data: data
                                            };
    endrule
endmodule
